`ifndef SONGPARA_VH
`define SONGPARA_VH

parameter song1={
    4'd0,4'd0, 4'd4, 4'd4, 4'd5, 4'd5, 4'd4, 4'd3,
    4'd3, 4'd2, 4'd2, 4'd1, 4'd1, 4'd0, 4'd4, 4'd4,
    4'd3, 4'd3, 4'd2, 4'd2, 4'd1, 4'd1, 4'd0, 4'd0
};
parameter song1len = 96;


parameter durations1 = {
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000
};
parameter durations1len = 192;

// "Mary Had a Little Lamb" with varied durations num=18
parameter song2 = {
    4'd2, 4'd1, 4'd0, 4'd1, 4'd2, 4'd2, 4'd2, 4'd1,
    4'd1, 4'd1, 4'd2, 4'd4, 4'd2, 4'd1, 4'd1, 4'd1,
    4'd2, 4'd2, 4'd2, 4'd1, 4'd2, 4'd1, 4'd0
};
parameter song2len = 92;

parameter durations2 = {
    25000000, 75000000, 25000000, 25000000, 25000000, 25000000, 75000000, 25000000,
    25000000, 75000000, 25000000, 75000000, 25000000, 25000000, 75000000, 25000000,
    25000000, 25000000, 25000000, 75000000, 25000000, 25000000, 75000000
};
parameter durations2len = 184;

// "Happy Birthday" melody num=19
parameter song3 = {
    4'd0, 4'd0, 4'd2, 4'd0, 4'd5, 4'd4,
    4'd0, 4'd0, 4'd2, 4'd0, 4'd7, 4'd5,
    4'd0, 4'd0, 4'd14, 4'd10, 4'd5, 4'd4,
    4'd7, 4'd9, 4'd10, 4'd5, 4'd7, 4'd4
};
parameter song3len = 96;

parameter durations3 = {
    50000000, 50000000, 50000000, 50000000, 50000000, 100000000,
    50000000, 50000000, 50000000, 50000000, 50000000, 100000000,
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    50000000, 50000000, 50000000, 50000000, 50000000, 100000000
};

parameter durations3len = 192;

// "Jingle Bells" chorus with varied durations num=20
parameter song4 = {
    4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd4, 4'd2, 4'd7, 4'd0, 4'd4,
    4'd9, 4'd9, 4'd9, 4'd9, 4'd9, 4'd7, 4'd7, 4'd7, 4'd7, 4'd7, 4'd4, 4'd4, 4'd4, 4'd2
};
parameter song4len = 92;

parameter durations4 = {
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    100000000, 50000000, 100000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    100000000
};
parameter durations4len = 200;

// "Ode to Joy" melody with varied durations num=21
parameter song5  = {
    4'd2, 4'd2, 4'd3, 4'd4, 4'd4, 4'd3, 4'd2, 4'd1, 4'd0, 4'd0,
    4'd1, 4'd2, 4'd2, 4'd1, 4'd1, 4'd2, 4'd4, 4'd3, 4'd2, 4'd1,
    4'd0, 4'd0, 4'd1, 4'd2, 4'd1, 4'd0
};
parameter song5len = 104;

parameter durations5 = {
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    50000000, 50000000, 50000000, 50000000, 75000000, 50000000, 50000000, 50000000,
    50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000, 50000000,
    75000000, 75000000
};

parameter durations5len = 208;

`endif