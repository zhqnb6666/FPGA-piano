module TopModule(
    input clk,  // Main clock
    input rst,  // Reset signal
    input [7:0] key_input,    // Key input for key.v
    input higher_8,           // Higher 8 bits of key_input
    input key_on,             // Key on signal from keyControl.v
    // Other global inputs like switches, buttons, etc.
    output [7:0] led_output,  // LED output from led.v
    output higher_8_led,      // Higher 8 bits of LED output
    output buzzer_output,     // Buzzer output from buzzer.v
    output [6:0] segment_output, // Segment output for display
    output [1:0] digit_select_output // Digit select output for display
    
);

// Inter-module signals
// wire [3:0] current_track;
wire [3:0] key_out;
wire [3:0] note_out;
wire key_out_on;
wire note_out_on;
wire [6:0] counter_value;
wire [6:0] time_in;
wire [6:0] time_out;
// assign counter_value = key_out;
assign time_in = counter_value;



// Instantiate keyControl module
keyControl keyControlModule(
    .clk(clk),
    .rst(rst),
    .key_on(key_on),
    .key(key_input),
    .higher_8(higher_8),
    .key_out(key_out),
    .key_out_on(key_out_on)
);

// Instantiate led module
ledControl ledModule(
    .clk(clk),
    .rst(rst),
    .current_track(note_out), // Connected from keyControlModule
    .playing(note_out_on),    // Connected from keyControlModule
    .led_output(led_output),
    .higher_8_led(higher_8_led)
);

PlaySong playSongModule(
    .clk(clk),
    .rst(rst),
    .key_on(note_out_on), // Connected from keyControlModule
    .key(note_out),      // Connected from keyControlModule
    .duration(counter_value)
);

timer timerModule(
    .clk(clk),
    .rst(rst),
    .time_on(key_on), // Connected from keyControlModule
    .time_in(time_in),
    .time_out(time_out)
);

// Instantiate buzzer module
buzzer buzzerModule(
    .clk(clk),
    .rst(rst),
    .key_on(note_out_on), // Connected from keyControlModule
    .key(note_out),       // Connected from keyControlModule
    .buzzer(buzzer_output)
);

// Instantiate DisplayCounter module
DisplayCounter displayCounterModule(
    .clk(clk),
    .rst(rst),
    .counter_value(time_out),
    .seg(segment_output),
    .digit_select(digit_select_output)
);


endmodule
